// module adder(
//   input  byte a, b,
//   output byte sum
// );
//   assign sum = a + b;
// endmodule

module dash();

struct person{
  reg a;
  reg b;
} person_t;

endmodule